PK   z��T@j��%  �A     cirkitFile.jsonśKo�6��J�^�@�z��m{�C���bC�$j#ԑ\YNv俗#'��R�� u�$"g�#��p(3�^��M�mg�{�m���Bͼ[ݕz\̼u�d}�}���֛?��_�h��mc�>+�rP��Ƣ�C����P�q�WJ�in�$���r�nuAS�����4uES���9eP��V��K!����ϣ ��*�*J󴌅�sB�1�e���к,%�J��H� J�J�Ii: 5M�f�8�DDԏ��D��z R�O�@��@����? �D��ȟ$�'/����G>׸IhZ�����:.ӄ�cJ˗VǤh��On�v�v����1^)�e�,V$���Ŋb�V
�U��h�JED+	��<�1��C���k�B���ߪ2* ���"�1��X�P<S�	�����b�x(���b�X�P,ߤ�5�������t@wM3��]הq����^����5f�wzEL��V�Ŋd��XQ,V"+1����J�C�<�
|��`�C��AX�0,x <���y(���b�x(���b�X�P,ߤ�9��[����	���X��_c���gY]~����{�;���+]�2��aە���7�P)9�rF� ���PZ&=�RӤG�[._��]{o!�My������'9@d�� �dR�ݕۺ�o!��mUy���.��ˌ����Q_�C��"�c���[�#k�ɐ�.��EƓ��g<�Q�Cyj��`A%x�9��TTL�S�r
�8J�@��@%�$�D��T�J���('Ht�ٹ8�-�[�u��-�Λ������^��%fi���4�!��'��_x��{�}+���'b�N�;E�A%�
�(,PZ��@y�
5 5`���������5�ppӥON���0�]?4��n�v��Nz�t���>��t���;>%�t䖸a>�ΤS����+K=>aY�ܬ�S���M�6w:�C�8���*8���U��^����7��vSf��U���M��8	�|�S凲�~����"�e
:Jt��?����d�2U��|��rO6��^۲ǡ�kצ�k3��u���g��������F}��X;���j�W?�=E8۷Mm��_����S���+��[�1ݗzS�+�/���ۺ3v�����q��m��~ۙnʁ��ȓݮ���е�����%7>�*V3��x Ul�]�h�l�+s4�?����~�K[b�2�{�;� >�ڮ��w�x۵-*�X��!���m&�`9Cw����jD<���5�F�kĨ&���Ԩ<�2�zP�۪�:��P���pJSNi�)�`BS$�"��TS�����*�\�L(�zjB/�Ѓ)G/�-���������//���+q��ϙ�t8+��FI���Y&�DB���W��3SY�"mChY�aag����/eE �0*?��N���̴s,LG�$��ֹs�Ip���|�To�#��)��޷6
z��`7��a��e�T�����oma����ޚ��-Jʑ�c���1}�ŭ)?엣�����/�y��_�2����O7�|�r�e��6�뮿����P��|n0f�rҔ[z7����gN׬�_��[�u�_��v���X,<\�?U�X�yXJ7X:����xQ��x�b����I���^h���g�=Q�b�#�-�ޓ�����1.N��Ę�D`%1����sd��ȳBveR����p�H̑�ݱDN��Q�(>�Gb19;��1�Ef���`�r�b��XNvFv$3;/;��Nzv�TQ�E�bHq[�V@L���S���MWۭ���,N���ǔ�ٝ�^}h�>��n�w�|��PK   ��T��N�5  �8  /   images/5277c62a-43df-4c39-a7ff-d396621a1e5b.png�{WTS[�.��bGD�)���Z�A�t�*R�$@l(�")
"H�tD1HR҂�P�B��8��<�3��>ݛX̙�����o+���f'�]8���s��Ԓ��`6��#���[�n�r4��=���L�����D�EC�M�0�ʸW��`��M��awDQ16[���0�L�y�jB�;[�pO�1� � �����|�a����~A�$�N���X��A��}=�լ_�G�Ux���W,�u�	��|N�.�w&8v���n	j��޷��-?kݖ5ί��7�kk���D��37#	����j��P2U�����D0�����;B���h���]4���,q4eҮg���V�!�����%!>�^�n�nJ}[�=�o=I͹v�į$���~X��������"���`z_<��sfu�����B;��+��x5�9V�'�!wDu�+d�`��'�}�j<Vw�6aQx��{�[��?u큍���e��"�z�5D���j*�����g����k���;x�,�T����D�p�j��!���ѿ�A��_�����D>�V&9�D�nd���5�4�n6[�Е}�1����YR��P�r���uR��t�� 2�M�7�0�^��7��s��RX���x啋�4R�W;^yо�o�����ᘿRitw3��@2���M�Z�(̖�O�`_��j}Z���OIuF�x�1�a��K����Z��%����-%�fY�
{�xq�О�'�ܕ��,��).Mg�}�e��/�;z��fds��׾�����נ�:�A*C��ԮJ����ӽ�8ǔ�rc��I"�[	�N�����:HvoB_l�_.�W��j������!28�U����5�՗��O|.�lB��N����7�j��I��T>;�{)���=&��ґ%h�.%b��e_��zr�����2΋*O�]iJ�@��^NX��ly2��E��n3�����������$�=���P97pnG)p�;�n���05Q����W����}���zэ�>��3��]��]���V�ӫ��|�e�) ��9��<�s�ݕ�����UeI�(�s�Cđ���ޟ&�R����z��Q�کw�}S��Ϭ<�:�5����nH;I�C+0��B5>FG�ٕ�Q�U��s�1��/�A��C3���}�,&����^��'�2�[7������,�i��Q�G���E6�7��ŵ�z<l�ݱ��3�ԈB�u�7����w rܮȸ��թD���h �6�v��l���`���BFlFEQ�ۡ�cO�;�[����+�&��0�ôE�2��n8"T�@�qH��46���A${f��91���$�������4�ϕ�F�Uo�����[��)8N�:�x�r��i��#W�H,_J�ii�|����}���e���\���i&�U���p�Qv��c۴7Llnbo��y�.]=������^'��X�<���IS�n�u�E��{�.�+Ѝ��̦�j�]��4���{�"���q1��i�Ҍ�4��d���u�֧��zVPP�;&������\;5��B�\S�^_��9~<�h���RJƐwg��iG�ۣ1S���Ҽ�s�؋"��MPO���88{����E��{ ��[�4}��8>���'%��qeh�2H�����~$����5���#�<5�L��:%�w���-H���;}�+t�����>�U`�e;-�ݸ�F�xs�L�=˧Dlr��(�����`*��i���#YK��gt�� �%��.l�����sER��U�3z�r}E��Lh��"�M��)�3*Ͷ�{��z�Й�Gkz���A�p�D��8;=]���q**�quAc�;"(�J��8Ȼ��y�}NR�3��i�{�+��bO�D�[��/������K���߬����ʠ5��G����%h�߿ߜU��m�˱t��_���#6���1=5������Ճ_K�������^�	�'.h�!�]�p�Y3n���MmO���()(�}�� �%1����R�t��D7�e1��/^�HHH�hdZ�_�v-W��(����W焌���l�R�P>I��C������ ��7u簒k��fDc���17��O5de�����6�q~���s[���-�6�@ǫ��B���%q[�C�)�4n�5�Ӎ�8���u{�$�S� ��px)jh��-�$]�����7�7�	�U��h1X�nOІs�I����>���P�_�F�3kw�x�^�_��@ɇ]�-3�^V6ֶM�8�B��ֵ��)��v��f���L5�3r�j��*+-#y������˓�΄��|*�>�iS6�9%��m�粩Q�4 ��Ƣ�-���gc��%N��q��N�V״�R�K����\^�z�?s�8�d��E{���B�C�]�<D��V�/�����#(��ڡ�&�?|�ŧ�u�#�[L��~�|�p����G{�H����@���H$0X����@3h��N���^j��c�ޞ����b��s��(���g
{'8�]������~N^y��[m<i��z�w@�����,��B.�X �`�������j;���#�bȔ%��yO�^�������kZ���[P��{���9UO���sW��,E\���4���$�-;�A}a{�D�b�t�ۿ�&WO� �e�K]@=���B�m_e>�9� ��u�� ���P;b`�϶�Q��*�%��+t�>E	���P�Z�����5"�T�����`˛ZW�m�:�t�Υ��ڢ���i����໓���m"#��PM><��_-}������kk�vp��P�BF����A�9�5ds��#}��%�C��m�f�����jM���@S;���=�/,���c�i���ρϒ`�7:�_Q�#~��>]<]��`�~��[ZrI��2t��
1��j�2�kRO���ӓ������ʲ�ZѰ�Դ�y��W2 �a�WdGQ����2�ޟ�V�^��T��)]s	)����朵��F�-�N.�5��+v!]�/Oz^���l��E)��,��PU` �-�qٓ�_����ggg���&��\��8�^�{�]깪�OX,���J���H�TXߔM{p�5�1�=+r
�.��?|p��U��YlA��p�=T򚁉t}R�Z7dΟ��'y,�/V�v�:�!�6B�{}z��^�'�VI܊hf�Y5m�*cukV"�ѫ�g�]E�f��E$�kX
U�I��y�3�{��os�@�Vm��c�ϓ)�-�<��*���꨾�v�2�s�wv=ԫ8�=-�#��4WV�\���#`A~Oz����?vM����ݗ;��ޕ��U�#�����V[��t"��a�[�Կ��֟PD�7{.Ja�&~��LL�l��0�rF�{�E����y:'�d$��q��ƀ��_��;$��T���;j��<�w%j��`��]=G�Z�J�%�=N��_���eM;�[ז�KJ�M������0֩,���@��Ֆ�y�x�9�3�#��]X�[���Ȳg=A�S�(J�t�Y�3�:�~�c�	=�`|ۙ�1f��;	�D;�U`/��L㼾y���u��9��.{Z�a��bX��s߻���wq��?���jm�]@��)�� շ{�轢�J��ҝ~�� �A���9p�^�Kc�����,�������+�kXe���`��$�Ɋ�6Y��MՙF���
�~��Lf����?�+����Z ӈ���s&4�!࿿�O��lm��k�{s[�n�xIc(�N>H��T����1]Cky�����[�%��D��D� �S�lU����X�h}�S�|]}��"��,��k������ϲɣ��)	�*��.\ko<�%`����L��x�=��x%��ۅ�u��j|�^镻�<��(���\j�3�L\�!jR�FB{��"��M\�Jz���=� 3��H�����7�+m�`�jM�x4�	�u�2�v�_w�dv=<}r�j�6R�߫*��ًsk�
��NS&�hѫ��^�gU�R�}����j�·CJБ�0�c*��J�mM�y-�,:4���S��E����U��qR/aK�Eg�V��c���?x������$5��
��+krz@LL=8F�2>�Ŋ�@��
����ɠ0,�bS���m?{-Y.AT�F�v�
(5��i�p%Z?�.�*�qPsz/bX�jt�)�t�TK}���'<�zM�����E�*���/��Bq���6�U���� �0|� %�wm�Ƅ>vڼz3M#��JrU���rm��Qڜ��z��������l�9%Qk?�	��***���d�	�xƄ�^��1/ߪT3��gϼ�������,K�Z|�j/`QjV�%��q�Y>*����Rȩ'U�oYg��5�D��J����(���.���ek�@����？���?.mV/�5���x$!Vb�ƈ5V���7��T=$Y��W���r5Wa|�OX�/�"��J6%g�I)��Ȇ[��@Q2lյ�M˭7-�%�ƚ�od3Y���ZV�9�.�ѥ�v`{����[���OZ���A�5>��3+B�N�4�ܕĝ��:c:���`��kKQg�ϋy~�2YY��av�Z�f��u�Y�ڞ�$��
�p��a,l�h�����=�[��ye�-�ާ�vYC4BƼ̡x
��'�M�md+яoU3d|]eNj2�
3�)�a	��3޲��	�n������Z�~"�a��L�V�4G�'f�p �<�Xb#�	Ҧk{z��� A����F�yw� Fˀ���XF�G�cY&��g��|1W�<LmirQ!��m}K���g2�z�����߲C>�+F�U�P_�(��]��ۜ��>=a�ۼB����*y�ϱo����3��3�b�a�̜�o$g�0N;0�G	r���g�� w��t�oS��'���1��9&�}�JI��iب�D��<g3�}�N�B�Q4co&�1>�0Yy:pc5�X��4�Q����>5e:)���,�DQ�|.�Ѓ��s�
-7��V�R�E���ג;�{:��Hߡ��z�_�������ξ�f��2�ͺ;�"\�*Nͮ�I��q	��>w4G6#�[R:����&¿*�
S|�=r�K>���?`\>J�=�5� �KeK0]�]ю��O����B�և�����-C}�Ӳ�P�0�xM�� R�í�-� �Sc�RӻE�C�ɲ��4�/�|MI���	k �:%��W����[|�Z?�֦����R5��!��|���18�3?��ᮦr	��hݘRJ�J�W<�^6^6�M��4Dn�|���w�5rP�i�U�,y9C��|C��\�O#^�3 �J���ZʌV��Yh�߅� 	ȼ��c�n~5�r-Ek�7^
��Ӗ2�R�(|\	�ַm��e����6wH̕H�'ᢌG�D� ����z��6f*�[��d�c������Q)uy�}�ჽ��t���m�c�.�[��u��"cQ1&^��o���a����T� ��:�5�b�`��AU;�}������0�(���D�G�
r��v�S���b��S0�k�LgJ��gAX�S
�uwP��`[�WD+J��K`w�>'�[҅Kab0Y-��!�*4Hǋ�8�K�£6r٤�t ��ĚX7#��%M�m�cZ$�z��4�z�ο����^*�2�Z�F���Q29�o73�"E��:����2�s��}�6J�h�S_��D�T,_@N�ͽ-�L������Y��$��� �܊��y �����	�a��(��ą���@��y 0����"6�u�dM�2�=t,2SG2�}� L&县j?e-5ͮ2�h/��ڮ*T%krgU�����m0���-�k��,Fte.��Y��W0Cko��$ݵ�@��T���n���k��m ��7z$��x�2!\m��"SUJ�ؐ�L�X���'�{���.-3���{���#��ᘔ��/$�|fH�xڋ�E5_fn�o�c:���z�2����U��0�
B� ��?�p�׻Z��MVQ��^���!�Y	Zy����Vɫ�eos&�,�}n�T�7�V�rF'w<���I�\&2��#k�5�������m1��7=4���q#�F!j��7���)�*�փ`�Hە�_���2���'� s����X�f�[}�7�}R1����/2�h?��J衴X��C�4*=s~
�������K�/�{C���iA�=����a�	F	Ao����Z�<\����*�u�s
YgB%|�v�b�	����<	�m�������{L�e�*�~�m��u|/��~��?Oy6��$)�S��ʊ���#��*���.^�5��ĵ4�H$�O&2��%�Wɨ���2���jt�%��͊�@B�:�s�Q�Eʍ[�G�������`�KqS?gD�<B��/�N|O��L���ߊ��Qs�4�@�lg������˙�Ԇ�q��_����������dU-u��+r��Sk)-yq�w0<Y�
f�$�.������*���5�3�62x�9T�VP�&!wd<w���-<���F��-nI�}�@�YI�q�s6{��M#fyO�J?㣛WQ��^�F8i3z(߿u���+��Ͼ	݉�Cm���{ުn;��>(s
�����}�������v�'��:��IiJ��! �J�{tn������q^���؈H2��l�6�."�a�qʖX�*eL]��h�Ϡ{R���s3�"�⚅�� �\�vM,"	���ڮ�z�2VD��̌	X3z� NDE�$�~4�{g���s��qZ)��6̣�mѫn��\t�S�XNzbω�a�h:}yЏ�Ȳ��f�oHd9��z��bI%�Z7�$������y�M���}LAoo7����=$5uY���� סH ��j�V�F�@�MI|kC?owF
�<�u��vj��ֳ��6�hR�s���eǀ���:��!]���^�iov���?�Xc��5��pVC��i�!�2f��aj�\>Qږ^G�A#�"O�n�Ι�q��ǕJ%������C5�l�:���=�C� �3/j�lǽ��~ ݱ���"��~6: ����[I�k������1��̄C���;�$w%Ε;I�&c�ZkڻOc�t�K�;ۦ��&�?�5w_3�#*(��h��w/���xx����;��6.ff⚯W*�qSc�CʞD(�ç�m����s�5��f�޹
�i� �ƖƏ�\�M��dz,�\�I��I� ����>��.���N�R���yX��YD�#�T�	̑;���^���Qas���.��z��F�q��罣~� m&�XnXN#bc̖��������Bn���/��&N���4�]z9vG�#�Y��^�<!'�j��0�vޱz�dMee�e�)���NR�Cޫ=vbsJ`����b�DqJ���L��4pʸv\;}Lx���ſe	��n��ᨄ�y^���?��չ��+X~/i�iw�%2Y�_�ᱍ(����n� \%�4\�k���{��|�)m)Ǽ]Sau�h��S�x5(���.3��Q"�.�@L���gy(� �7o`U� ��G޵��R.u�NT���_�f_&r���lNg~�r�q��G�H�;<QE:N3�/����$�v�,c���9�kjL1o&���!F����Xm��<O�����#�d���������ė���>��4�-^�t���8 �'��z}�A�|���C{�i\��t�)e��H=�ֆ�����ORN����?���T^�%��	��Q��re��D�� v����Mc��y��G10��+��p��"VF��/ÒL&�����'��`=
m����i�����$�Ӏ[�	������\�A��k6��G��d��q�/����?9)�[�?,Ӣ5Z~>m!�J����7}�(k�
diN[5&��Y��6�j� �Nc��4�cL��N��$ j3o��v�S���.�O��w_<����Ax��;Yh��`�����3�{"�3҄�A�8(���&�&{e��^�OII�W��O�M�SMQ%R]�?Q٣$�2(�%�-Ԝ�#ݒ��� �ć��'1�*T����'�Е�� � ��?}.zօ�"���qF'VRb��
.J��O͑?��#+e`��,S|�飒�\���\�S(��U��Lr����i_v�ѕ^l��/��r�?�������d�Y}��L�H_{%7��8���ß�z�bă����`�T��#�f�� �j^��J�+7L��㷟����w�S��<kdo���C��lJj����G��r�S�X3��� 4���S>
��k}�����?LÔ�h�H�ۯ���9+�r7���$8�
)>.�vւT�l�� ���A����^$�����]w������'$H�$��6{c��a��|�&߸!�4J�����?5�?��R���a�N�i�˻�A/9���C��Y'�R ��1�?'0cP�L- h�d�z{gR?�2��y6n� ���e`�E���f�S,���uR��SRM�����6M�%C�Vz��v�<_��cI�@cpd��kˎ���n�����b9`�^�Q������Z@ٜO�݆���%
���K����&�L5�������M��Sry}+���xj���}+�������le	X�KW��hcG��W�������G\����8����?����_4��U��ڣ8ڹ򶟮7<X��Yf6���L��&�ɯL����q^u'yJ��1����~jC�Sv7;O2�5x:.]�}���6Zoi���Kp�1,�HU�!Z/�W��R����up��|�_x�о_w��6�M&�q���î,[��� M�K�z�k�7��[���˼9Ee @AV�����	��Y�Z8n�*�o9����)��N�a�9�-�cbVmͧ����#t�&ܾvI�L^>X{�rΣ��~HziH����va�yU�Pt�6�d���Hc��g��Q˯���u��)�����ozz�_)�.W���$QV��:�\3OT�L�j�a����܄�|W�O�^ϓ�ъ�1���:7�̸�P��fIV���@������rX���T���@s�F�9m�0�!W
4�
7�6�CțzE�+A�wcq\�m������rObGߟ#�^�g+ЇT���s��.��fį<$[�%�y�����۽΄J�
����6��Z�.V� ��L��*�: ޢ��/m�UH@�lp|i�G<_V���K�������!�?��:Z��;h�^��wP��=ر�f)����̊7�F���a@��8S�<�mN�ѿ}�M��� 9m���ip�z"�7�/�zP/ZrЂ��rl���v�b�����R"�f.���yֻ����W�\��I� ���_	��n�w:A��J �Ƹ���w����� u{��'@��c�5?��	�o�,���n�Ư<7{#༗#��
�}�^�|������'�?�͞7��������ǂG��{o�����w��AC��?0�M��S�Ck?����GC�y+,Ĺ�������Տ��$fM����������|?4}˶֬��t0�7A޵����1��4^XC�*�+���H�=I
taz��~��,��u�@����Uer���y���2d��$�?G�+��wT!%F��܁w��Vs��x�ۍ��L�W�gi�<��F�����}�w�?��}Á��W�%��Ue@֩��#����g�����ņ2E�v���%��N�s}`��6��4��Q`�>Ś����|��>Ǳ�*��>���n}5�'&�`��J��W�U�DpoQor�[<��q��3�6��3w�����S�����֗J�;�b̂�`��(�FËm·���2��K�7T��]����������$GаU����>��W�af���?�C�U�o�U�$�G��~��%�0*����b�&�Ѓb�.H �C3��ƶ7�,�jD���!8�cS�~Ot h�(�&.e�m�Z�ї�E��2�i���h�ӭ/oM u�Y�#����d+;�f�c90�rwBȍ�R�l����Pz�A��s�����̥T�>l�mA7Y6��p|���Jh�~�S�<<w_�>}~�ޑK}��>AL�ݼ!��%:§�i��� ���Dp�_����/R�|`ڂL��#�lݪ�7��Q!��/8�L/���h��<a�hQ������k���cp�^��2��18�[�`�x~=!7��-���d�A��|�Eb0z0�㲴&��K��M���j@�f��?d�"o|3s�܊�*�:�/�0i`D6�}GTt���]��8 f��z�C*O�A�1��2�4Q 7ΰ���^|'�B��έ@�f�~���l"G/���P�B�F��I n?H��靳�rY�q�+�)��%�k�T���l����m+���C% K�2ɁU�����@.�,�?����&�~ۃh�M�I������n�#Y�� ��q�&6F����s)'������Ml�d�����t���c�M�����@(�x�_�nb�p ������p��@m��+���@�j�Q^Tz�2΀���tw�jiiY^^�R ͘�o|��4�Y�)D�Fk��Z^p˹���րI�>��ͼ9j,�0>��X�K��G���S��<aַ�w?:������l���Vٔ��-/`��3�bNV�* S�8G�!��+?�˹�.C��a�7k�e��N�X����yg�-���;���%:����&oM�|!5�H��=�}�4�Yq��I^2�,�Ay�t���,�o� Ҍ���5���O�ִA���j�\�/T��@fVVUIDQW�_��A�-?$t�وf��`g��U@}f��[s�C.�}z����M�R�"�WA���n�A�D!����χ}޶"xb���|w��7���s�����N���Q����ֽ���$�tYڇLn��u����]Gs�@@g_�f�i��ϓ�������_w}oAe��ܨ��i�t�����R9����E�vT���è�&���A/[����_J߇2�R���6���.�����.�;}��j�+����ng�:��~�#QôsX��EV��7PF��^���X�:^����6v�\1w�&��0�������B&�%@RbIoE��&D���v.%���.�2<�4[|y���g��/�Q����=S$>=�L�pHs��3җ�ӄ�+�{��!t|�6���Q�+?��]�	�]K�z��;�G�}uUH�鷂�.��S�\���W��滐*ӓ�n�&�c}��ϊ�S8��}1�^w�;��FS����W&��<HKP���8�;{+����Y� �G�F�B<��_�H��Ο�|�������g~�q����3��������m�T�2��'w� %v���G�Tgz�{�g'��.X�!z�K#��A	����r����׽%|�ovd��߿����@'A����|�:�W��VCm\�����Ėw����iL��5�� ��X�(�|G����W"r�G��M�ܸ����쯟���ϵ)�G�	��];٨�իԃ�.uN���%�����Жˉ���J��� �~�cR.8��+RkNYg
���*��k���b���L����f�]��-�"�������j(k�(g%`�������ŕ�����$(5	G��fqY1weҨ��ᲅc8ccQ�0�� 8s(n�3���PR\|���ȝ��e���?� ,�6V��+Ŏ����)o[(�D�666.**ҋ�d+e�~i:��S�ӕ�ץ�9����·6��:;;}||0��$<�&�s������i%E���Zޭa�HwTnotN�!��������e	r=>h3��>��0�L�f�S��~L���?�Q�wZ��}K����ue�����4$42�UU�[��qV�{u�$W��璼璏[�g�X"l�ٯ!�{��PfS&��?H�6���U�|��l�32CՅ�DF55n�1.�_�Z*�y��!���d;;;�mtĦ����!�BV�l��y��@������ӻ�"V��P1�a-�"k<ignn��[GG���C�'k�<~�_6�'��bOY7�.��uUrfF��M8�׮o��-P������`�q���Ǉ� @�.��~��u�����Yf�Y�����	�h��ౝ����0_�jn?� ����{�H]	ee�è�Q[������~���L��Ս��I @Z:�EC(8\�dñ��G?�TF�>\�o�WVZ*Bo�(��<XF{~���V��<���I�=�6�V���M����&s���5m�����c;Xs�NC���} ��%�Ѓ\#%2/�/BN��/�S�[���0�)�?�:tms�@�-U	S��گa-�ƴ�Y�M�$2�h"��ܤ���bI���X 9�FN� ǩ�K*!�)��`�����#�nV�׌���� R���L7���|���41�T��'YY^��ؘ���O�6[���ΨФ��y��d;��G|"�h�d��>�si�ռIl+7D�E׃n�/��D��ُ�#���b{����[�$��h���J�q�����@ԋi����+����;s>�� Bs�6a���_iE9c����E�-F�<�ZX�K�+�m�~��Pzl��3�'s����H ��yԐ���ĻrM�n��<e5��Rkz|w=R�0�ww��[O�,�ƒx���JVV0��A���z��h���1�����QC��.p�!ĭ8���߀��S��	��=%GH��B�f�������
R�z��:a��1���ݾ�(�`��1�b��%�ԽL�F;��ҭ� �b�[ڴB��4��T�,����4X��������{HHGp!�=�x�z��ZS�l�d��?C�!�~%p�p�:r��$���m��k"��Eg1CE�T!O�&��6D]�P�^��E����9�"�f�&�@(�x��R�a�wl��%��{>�i��~��HvݹZGC�j��^u�7��yB��QQѿ���=����%Mu�S�==������*�u���$@������������G'!���tAA\2�r���R�'L��qz�NOx1ʲ�Ɏ���r�F�J���@
���:����sf&��kk4G}7�Ux�s�@\�N^���zNk��:"e�~�����_��\a�k��)��ko���q�aן$�@��b}�^�ol��|H�8��O��j&�1�6y�`az�{�v�g���	���SЎ�7:zI�9��S#�7���D�Y�+_ju�cƢ��8�� �v{Gj)*�����\�u�z��imR�B����9��`��y�e���p���b�y]�����yio���ew'}nC�C��@$!��i�U����pI���	���'�f�JQ���"&�)6��\��O���F5e@l��f�R����PK   z��TNe�=       jsons/user_defined.json���n�0�_%�؀����Ъ�ϩ�*ǘt%bSE��uh�K��z�;�1��鎭"%靲o��A���SYF� ��(��o�ԑ��t��{�*��6):�3��"���꛸	T(�(�2�"LYU��dE(x]�+�&"Q�9>��Zv�W?�_)'-�����L|���Z�k]R����+pm#����	-�8�
��u�h~����l�������#�u��Y@>�����O�C���򈧜�(w�廱h�lڈ��z2���it:��E���4;[��ͦ�|v�����ck`�!>Y�*�����l��?Vb�_PK
   z��T@j��%  �A                   cirkitFile.jsonPK
   ��T��N�5  �8  /             R  images/5277c62a-43df-4c39-a7ff-d396621a1e5b.pngPK
   z��TNe�=                 �<  jsons/user_defined.jsonPK      �   ->    